module LedBlinker (
	i_clk
	i_en
	i_switch_1
	i_switch_2
	o_led
);

parameter

//1 HZ enable generator
always @(posedge clk)
begin
end


//Lit up the LED when enabled

endmodule