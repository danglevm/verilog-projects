module HALF_ADDER (
	i_INPUT
	o_CARRY_OUT,
	o_SUM
);