module ALU (

);