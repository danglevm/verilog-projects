module FULL_ADDER_4_BIT (
	i_FOUR_A,
	i_FOUR_B,
	o_4BIT_SUM,
	o_CARRY_OUT
);

input [3:0] i_FOUR_A;
input [3:0] i_FOUR_B;
output [3:0] o_4BIT_SUM;
output o_CARRY_OUT;

endmodule 